`ifndef ACCUM_REF_MODEL_PKG
`define ACCUM_REF_MODEL_PKG

package accum_ref_model_pkg;

   import uvm_pkg::*;
   `include "uvm_macros.svh"

   import accum_agent_pkg::*;

  `include "accum_ref_model.sv"
endpackage

`endif



