`ifndef ACCUM_SEQ_LIST 
`define ACCUM_SEQ_LIST

package accum_seq_list;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import accum_agent_pkg::*;
	import accum_ref_model_pkg::*;
	import accum_env_pkg::*;
	
	`include "accum_basic_seq.sv"
endpackage

`endif
