`ifndef ACCUM_TEST_LIST 
`define ACCUM_TEST_LIST

package accum_test_list;
	import uvm_pkg::*;
	`include "uvm_macros.svh"
	
	import accum_env_pkg::*;
	import accum_seq_list::*;
	
	`include "accum_basic_test.sv"
endpackage 

`endif





